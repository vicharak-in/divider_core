`define TOTAL_APPS 2

`define DIVIDER_UNSIGNED 1
`define DIVIDER_SIGNED 2

`define VERSION "1.2.1"

`define GET_DATA_RAH(a) rd_data[a * RAH_PACKET_WIDTH +: RAH_PACKET_WIDTH]
`define SET_DATA_RAH(a) wr_data[a * RAH_PACKET_WIDTH +: RAH_PACKET_WIDTH]
